CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
10
7 Pulser~
4 55 179 0 10 12
0 11 12 4 13 0 0 5 5 2
7
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
8585 0 0
2
41828.5 0
0
6 74112~
219 328 197 0 7 32
0 3 3 4 3 3 6 7
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 1 0
1 U
8809 0 0
2
5.89668e-315 0
0
14 Logic Display~
6 426 161 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5993 0 0
2
5.89668e-315 0
0
14 Logic Display~
6 395 143 0 1 2
12 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8654 0 0
2
5.89668e-315 0
0
7 Ground~
168 118 291 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7223 0 0
2
5.89668e-315 0
0
12 SPDT Switch~
164 263 101 0 10 11
0 3 3 2 0 0 0 0 0 0
1
0
0 0 4720 0
0
3 SET
-12 -15 9 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
3641 0 0
2
5.89668e-315 5.3568e-315
0
12 SPDT Switch~
164 200 135 0 10 11
0 3 3 2 0 0 0 0 0 0
1
0
0 0 4720 0
0
1 J
-4 -15 3 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
3104 0 0
2
5.89668e-315 5.34643e-315
0
12 SPDT Switch~
164 200 206 0 10 11
0 3 3 2 0 0 0 0 0 0
1
0
0 0 4720 0
0
1 K
-4 -15 3 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
3296 0 0
2
5.89668e-315 5.30499e-315
0
12 SPDT Switch~
164 263 240 0 10 11
0 3 3 2 0 0 0 0 0 0
1
0
0 0 4720 0
0
5 RESET
-17 -15 18 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
8534 0 0
2
5.89668e-315 5.26354e-315
0
2 +V
167 148 49 0 1 3
0 3
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
949 0 0
2
5.89668e-315 0
0
18
5 0 3 0 0 0 0 2 0 0 14 2
328 209
328 209
3 0 4 0 0 0 0 2 0 0 18 2
298 170
298 170
1 0 3 0 0 0 5 2 0 0 15 2
328 134
328 134
1 6 6 0 0 4224 0 3 2 0 0 2
426 179
358 179
1 7 7 0 0 4224 0 4 2 0 0 2
395 161
352 161
3 0 2 0 0 4096 0 7 0 0 9 2
183 139
118 139
3 0 2 0 0 0 0 8 0 0 9 2
183 210
118 210
3 0 2 0 0 4096 0 9 0 0 9 2
246 244
118 244
3 1 2 0 0 8320 0 6 5 0 0 3
246 105
118 105
118 285
2 0 3 0 0 4096 8 6 0 0 13 2
246 97
148 97
2 0 3 0 0 0 8 7 0 0 13 2
183 131
148 131
2 0 3 0 0 0 8 8 0 0 13 2
183 202
148 202
1 2 3 0 0 4224 8 10 9 0 0 3
148 58
148 236
246 236
1 0 3 0 0 4224 0 9 0 0 0 3
280 240
328 240
328 203
1 0 3 0 0 4224 5 6 0 0 0 3
280 101
328 101
328 140
1 4 3 0 0 4224 9 8 2 0 0 4
217 206
289 206
289 179
304 179
1 2 3 0 0 4224 10 7 2 0 0 4
217 135
289 135
289 161
304 161
3 0 4 0 0 4224 0 1 0 0 0 2
79 170
304 170
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
196938 1079360 100 100 0 0
0 0 0 0
1 66 162 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 2 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
