CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
17
7 Pulser~
4 89 239 0 10 12
0 15 16 3 17 0 0 5 5 4
8
0
0 0 4656 0
0
2 V4
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
9342 0 0
2
41828.5 0
0
2 +V
167 510 481 0 1 3
0 5
0
0 0 54256 692
2 5V
7 -2 21 6
2 V3
7 -12 21 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3623 0 0
2
5.89668e-315 0
0
2 +V
167 510 384 0 1 3
0 6
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3722 0 0
2
5.89668e-315 0
0
7 Ground~
168 85 138 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8993 0 0
2
5.89668e-315 0
0
2 +V
167 86 42 0 1 3
0 4
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3723 0 0
2
5.89668e-315 0
0
14 Logic Display~
6 197 59 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6244 0 0
2
5.89668e-315 0
0
14 Logic Display~
6 605 419 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6421 0 0
2
5.89668e-315 0
0
14 Logic Display~
6 582 401 0 1 2
12 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7743 0 0
2
5.89668e-315 0
0
5 7474~
219 510 455 0 6 22
0 6 4 3 5 9 10
0
0 0 4720 0
4 7474
7 -60 35 -52
3 U4A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 0 2 1 4 0
1 U
9840 0 0
2
5.89668e-315 0
0
12 SPDT Switch~
164 138 100 0 10 11
0 4 4 2 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
6910 0 0
2
5.89668e-315 0
0
14 Logic Display~
6 597 260 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
449 0 0
2
5.89668e-315 0
0
14 Logic Display~
6 595 150 0 1 2
12 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8761 0 0
2
5.89668e-315 0
0
9 Inverter~
13 239 296 0 2 22
0 4 8
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
6748 0 0
2
5.89668e-315 0
0
10 2-In NAND~
219 480 278 0 3 22
0 12 13 11
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
7393 0 0
2
5.89668e-315 0
0
10 2-In NAND~
219 480 168 0 3 22
0 14 11 12
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
7699 0 0
2
5.89668e-315 0
0
10 2-In NAND~
219 336 287 0 3 22
0 3 8 13
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
6638 0 0
2
5.89668e-315 0
0
10 2-In NAND~
219 337 159 0 3 22
0 4 3 14
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
4595 0 0
2
5.89668e-315 0
0
20
0 3 3 0 0 8320 0 0 9 11 0 3
153 230
153 437
486 437
1 0 4 0 0 4096 0 17 0 0 9 2
313 150
197 150
1 4 5 0 0 4224 0 2 9 0 0 2
510 466
510 467
1 1 6 0 0 4224 0 3 9 0 0 2
510 393
510 392
0 2 4 0 0 8320 0 0 9 9 0 3
197 296
197 419
486 419
3 1 2 0 0 4224 0 10 4 0 0 3
121 104
85 104
85 132
2 1 4 0 0 8320 7 10 5 0 0 3
121 96
86 96
86 51
1 0 4 0 0 0 0 10 0 0 9 2
155 100
197 100
1 1 4 0 0 0 0 6 13 0 0 3
197 77
197 296
224 296
0 1 3 0 0 0 0 0 16 11 0 3
271 228
271 278
312 278
2 3 3 0 0 128 0 17 1 0 0 4
313 168
271 168
271 230
113 230
2 2 8 0 0 4224 0 13 16 0 0 2
260 296
312 296
1 5 9 0 0 4224 0 7 9 0 0 2
605 437
540 437
1 6 10 0 0 4224 0 8 9 0 0 2
582 419
534 419
2 0 11 0 0 12416 0 15 0 0 17 5
456 177
438 177
438 192
554 192
554 278
0 1 12 0 0 8320 0 0 14 18 0 5
539 168
539 241
436 241
436 269
456 269
3 1 11 0 0 0 0 14 11 0 0 2
507 278
597 278
3 1 12 0 0 0 0 15 12 0 0 2
507 168
595 168
3 2 13 0 0 4224 0 16 14 0 0 2
363 287
456 287
3 1 14 0 0 4224 0 17 15 0 0 2
364 159
456 159
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
196938 1079360 100 100 0 0
0 0 0 0
1 66 162 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 2 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
