CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
100 510 1 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
177209362 0
0
6 Title:
5 Name:
0
0
0
25
13 Logic Switch~
5 810 800 0 1 11
0 3
0
0 0 21360 512
2 0V
-7 -16 7 -8
2 K2
-7 -25 7 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3221 0 0
2
41828.5 0
0
13 Logic Switch~
5 827 614 0 1 11
0 18
0
0 0 21360 512
2 0V
-7 -16 7 -8
2 J2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3215 0 0
2
41828.5 1
0
13 Logic Switch~
5 545 620 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
7 PRESET2
-24 -26 25 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7903 0 0
2
41828.5 2
0
13 Logic Switch~
5 548 660 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
6 CLEAR2
-21 -26 21 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7121 0 0
2
41828.5 3
0
13 Logic Switch~
5 291 668 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
6 PRESET
-20 -26 22 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4484 0 0
2
41828.5 4
0
13 Logic Switch~
5 232 685 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
5 CLEAR
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5996 0 0
2
41828.5 5
0
13 Logic Switch~
5 289 727 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 J
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7804 0 0
2
41828.5 6
0
13 Logic Switch~
5 230 757 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 K
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5523 0 0
2
41828.5 7
0
13 Logic Switch~
5 476 431 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 K
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3330 0 0
2
41828.5 8
0
13 Logic Switch~
5 474 332 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 J
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3465 0 0
2
41828.5 9
0
9 Inverter~
13 752 763 0 2 22
0 3 17
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U4B
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
8396 0 0
2
41828.5 0
0
9 Inverter~
13 270 757 0 2 22
0 8 5
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
3685 0 0
2
41828.5 0
0
7 74LS109
18 424 703 0 14 29
0 2 11 10 9 5 7 6 2 15
14 16 4 12 13
0
0 0 13040 0
7 74LS109
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
133 %D [%16bi %8bi %1i %2i %3i %4i %5i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %8o %9o %10o %11o %12o %6o %7o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 5 1 2 3 6 7 12 11
15 14 13 10 9 4 5 1 2 3
6 7 12 11 15 14 13 10 9 0
65 0 0 0 1 0 0 0
1 U
7849 0 0
2
41828.5 10
0
7 Pulser~
4 337 586 0 10 12
0 25 26 2 27 0 0 5 5 2
8
0
0 0 4656 0
0
2 V5
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
6343 0 0
2
41828.5 11
0
9 2-In AND~
219 676 747 0 3 22
0 17 12 4
0
0 0 624 512
6 74LS08
-21 -24 21 -16
3 U5A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
7376 0 0
2
41828.5 12
0
9 2-In AND~
219 680 655 0 3 22
0 13 18 16
0
0 0 624 512
6 74LS08
-21 -24 21 -16
3 U5B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
9156 0 0
2
41828.5 13
0
14 Logic Display~
6 560 802 0 1 2
12 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Q2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5776 0 0
2
41828.5 14
0
14 Logic Display~
6 588 811 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 Qn2
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7207 0 0
2
41828.5 15
0
14 Logic Display~
6 329 795 0 1 2
12 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Q1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4459 0 0
2
41828.5 16
0
14 Logic Display~
6 380 798 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 Qn1
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3760 0 0
2
41828.5 17
0
14 Logic Display~
6 748 328 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Qn
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
754 0 0
2
41828.5 18
0
14 Logic Display~
6 709 329 0 1 2
12 20
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 Q
-5 -22 2 -14
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9767 0 0
2
41828.5 19
0
9 2-In AND~
219 524 323 0 3 22
0 19 22 24
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
7978 0 0
2
41828.5 20
0
9 2-In AND~
219 524 440 0 3 22
0 21 20 23
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3142 0 0
2
41828.5 21
0
13 SR Flip-Flop~
219 624 406 0 4 9
0 24 23 19 20
0
0 0 4720 0
4 SRFF
-14 -53 14 -45
2 U1
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
3284 0 0
2
41828.5 22
0
28
3 8 2 0 0 4224 0 14 13 0 0 4
361 577
470 577
470 667
456 667
3 1 2 0 0 16 0 14 13 0 0 4
361 577
381 577
381 667
392 667
1 1 3 0 0 8320 0 11 1 0 0 3
755 781
755 800
798 800
12 3 4 0 0 4224 0 13 15 0 0 4
462 703
644 703
644 747
651 747
2 5 5 0 0 4224 0 12 13 0 0 4
291 757
370 757
370 703
386 703
7 1 6 0 0 8320 0 13 20 0 0 5
386 739
348 739
348 824
380 824
380 816
6 1 7 0 0 8320 0 13 19 0 0 5
392 730
310 730
310 826
329 826
329 813
1 1 8 0 0 4224 0 8 12 0 0 2
242 757
255 757
1 4 9 0 0 8320 0 7 13 0 0 5
301 727
301 711
360 711
360 694
392 694
1 3 10 0 0 4224 0 6 13 0 0 2
244 685
386 685
1 2 11 0 0 4224 0 5 13 0 0 4
303 668
361 668
361 676
386 676
0 2 12 0 0 8320 0 0 15 17 0 5
547 730
547 771
705 771
705 756
696 756
1 0 13 0 0 12416 0 16 0 0 16 5
700 646
719 646
719 715
575 715
575 739
10 1 14 0 0 4224 0 13 4 0 0 4
462 685
528 685
528 660
536 660
9 1 15 0 0 8320 0 13 3 0 0 4
462 676
516 676
516 620
533 620
14 1 13 0 0 0 0 13 18 0 0 5
462 739
575 739
575 837
588 837
588 829
13 1 12 0 0 0 0 13 17 0 0 5
456 730
547 730
547 828
560 828
560 820
11 3 16 0 0 4224 0 13 16 0 0 4
456 694
648 694
648 655
655 655
1 2 17 0 0 4224 0 15 11 0 0 3
696 738
755 738
755 745
1 2 18 0 0 4224 0 2 16 0 0 4
815 614
737 614
737 664
700 664
0 1 19 0 0 4096 0 0 21 24 0 3
678 388
748 388
748 346
0 1 20 0 0 4096 0 0 22 23 0 3
670 370
709 370
709 347
4 2 20 0 0 12416 0 25 24 0 0 6
648 370
670 370
670 470
492 470
492 449
500 449
3 1 19 0 0 12416 0 25 23 0 0 6
654 388
678 388
678 270
494 270
494 314
500 314
1 1 21 0 0 4224 0 9 24 0 0 2
488 431
500 431
1 2 22 0 0 4224 0 10 23 0 0 2
486 332
500 332
3 2 23 0 0 8320 0 24 25 0 0 4
545 440
592 440
592 388
600 388
3 1 24 0 0 4224 0 23 25 0 0 4
545 323
592 323
592 370
600 370
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
196938 1079360 100 100 0 0
0 0 0 0
1 66 162 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 2 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
