CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
8
13 Logic Switch~
5 117 156 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -15 8 -7
1 T
-3 -25 4 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9466 0 0
2
41828.5 0
0
13 Logic Switch~
5 120 119 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
5 CLEAR
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3266 0 0
2
41828.5 0
0
13 Logic Switch~
5 167 110 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
6 PRESET
-20 -26 22 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7693 0 0
2
41828.5 0
0
14 Logic Display~
6 168 210 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3723 0 0
2
41828.5 0
0
14 Logic Display~
6 198 210 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3440 0 0
2
41828.5 0
0
9 Inverter~
13 174 156 0 2 22
0 5 4
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
6263 0 0
2
41828.5 0
0
7 Pulser~
4 103 49 0 10 12
0 9 10 8 11 0 0 5 5 4
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
4900 0 0
2
5.89668e-315 0
0
7 74LS109
18 253 137 0 14 29
0 8 7 6 5 4 2 3 12 13
14 15 16 17 18
0
0 0 4848 0
7 74LS109
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
133 %D [%16bi %8bi %1i %2i %3i %4i %5i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %8o %9o %10o %11o %12o %6o %7o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 5 1 2 3 6 7 12 11
15 14 13 10 9 4 5 1 2 3
6 7 12 11 15 14 13 10 9 0
65 0 0 512 1 0 0 0
1 U
8783 0 0
2
5.89668e-315 0
0
8
6 1 2 0 0 8336 0 8 4 0 0 5
221 164
184 164
184 236
168 236
168 228
7 1 3 0 0 8320 0 8 5 0 0 5
215 173
211 173
211 236
198 236
198 228
2 5 4 0 0 8320 0 6 8 0 0 4
195 156
203 156
203 137
215 137
0 1 5 0 0 4096 0 0 6 5 0 2
141 156
159 156
1 4 5 0 0 12416 0 1 8 0 0 4
129 156
141 156
141 128
221 128
1 3 6 0 0 4224 0 2 8 0 0 2
132 119
215 119
1 2 7 0 0 4224 0 3 8 0 0 2
179 110
215 110
3 1 8 0 0 4224 0 7 8 0 0 4
127 40
207 40
207 101
221 101
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
196938 1079360 100 100 0 0
0 0 0 0
1 66 162 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 2 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
