CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
15
13 Logic Switch~
5 85 369 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 D
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8885 0 0
2
41828.5 0
0
13 Logic Switch~
5 145 335 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
6 PRESET
-20 -26 22 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3780 0 0
2
41828.5 0
0
13 Logic Switch~
5 145 417 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 8 8 16
5 CLEAR
-16 21 19 29
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9265 0 0
2
41828.5 0
0
13 Logic Switch~
5 123 113 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 D
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9442 0 0
2
5.89668e-315 0
0
14 Logic Display~
6 267 369 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Qn
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9424 0 0
2
41828.5 0
0
14 Logic Display~
6 239 351 0 1 2
12 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 Q
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9968 0 0
2
41828.5 0
0
5 4013~
219 157 405 0 6 22
0 4 2 3 5 6 7
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U3A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 0 2 1 3 0
1 U
9281 0 0
2
41828.5 0
0
7 Pulser~
4 57 176 0 10 12
0 15 16 8 3 0 0 5 5 5
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
8464 0 0
2
5.89668e-315 0
0
9 Inverter~
13 160 224 0 2 22
0 10 9
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U2A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
7168 0 0
2
5.89668e-315 0
0
14 Logic Display~
6 524 218 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Qn
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3171 0 0
2
5.89668e-315 0
0
14 Logic Display~
6 524 113 0 1 2
12 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 Q
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4139 0 0
2
5.89668e-315 0
0
10 2-In NAND~
219 395 236 0 3 22
0 12 14 11
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
6435 0 0
2
5.89668e-315 0
0
10 2-In NAND~
219 395 131 0 3 22
0 13 11 12
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
5283 0 0
2
5.89668e-315 0
0
10 2-In NAND~
219 241 245 0 3 22
0 8 9 14
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
6874 0 0
2
5.89668e-315 0
0
10 2-In NAND~
219 241 122 0 3 22
0 10 8 13
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
5305 0 0
2
5.89668e-315 0
0
17
1 2 2 0 0 4224 0 1 7 0 0 2
97 369
133 369
4 3 3 0 0 8320 0 8 7 0 0 4
87 176
114 176
114 387
133 387
1 1 4 0 0 4224 0 2 7 0 0 2
157 335
157 348
1 4 5 0 0 4224 0 3 7 0 0 2
157 417
157 411
1 5 6 0 0 4224 0 5 7 0 0 2
267 387
187 387
1 6 7 0 0 4224 0 6 7 0 0 2
239 369
181 369
0 1 8 0 0 4096 0 0 14 8 0 3
204 165
204 236
217 236
2 3 8 0 0 12416 0 15 8 0 0 4
217 131
204 131
204 167
81 167
2 2 9 0 0 8320 0 9 14 0 0 3
163 242
163 254
217 254
0 1 10 0 0 4224 0 0 9 11 0 2
163 113
163 206
1 1 10 0 0 0 0 4 15 0 0 2
135 113
217 113
0 2 11 0 0 8192 0 0 13 14 0 5
448 236
448 159
354 159
354 140
371 140
0 1 12 0 0 8320 0 0 12 15 0 5
459 131
459 203
354 203
354 227
371 227
1 3 11 0 0 4224 0 10 12 0 0 2
524 236
422 236
1 3 12 0 0 0 0 11 13 0 0 2
524 131
422 131
3 1 13 0 0 4224 0 15 13 0 0 2
268 122
371 122
3 2 14 0 0 4224 0 14 12 0 0 2
268 245
371 245
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
