CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
9
7 Pulser~
4 283 232 0 10 12
0 10 11 3 12 0 0 5 5 5
7
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3187 0 0
2
41828.5 0
0
14 Logic Display~
6 569 194 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
762 0 0
2
41828.5 0
0
14 Logic Display~
6 541 174 0 1 2
12 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
39 0 0
2
41828.5 0
0
2 +V
167 226 74 0 1 3
0 6
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9450 0 0
2
41828.5 0
0
7 Ground~
168 201 350 0 1 3
0 9
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3236 0 0
2
41828.5 0
0
5 4027~
219 457 230 0 7 32
0 9 6 3 6 9 4 5
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U1A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 1 0
1 U
3321 0 0
2
41828.5 0
0
12 SPDT Switch~
164 362 296 0 3 11
0 9 6 9
0
0 0 4720 0
0
2 S4
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
8879 0 0
2
41828.5 0
0
12 SPDT Switch~
164 270 178 0 10 11
0 6 6 9 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 S2
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
5433 0 0
2
41828.5 0
0
12 SPDT Switch~
164 361 119 0 3 11
0 9 6 9
0
0 0 4720 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
3679 0 0
2
41828.5 0
0
13
3 3 3 0 0 4224 0 6 1 0 0 4
433 203
333 203
333 223
307 223
6 1 4 0 0 4240 0 6 2 0 0 2
487 212
569 212
7 1 5 0 0 4224 0 6 3 0 0 3
481 194
541 194
541 192
0 4 6 0 0 8192 0 0 6 5 0 3
368 193
368 212
433 212
1 2 6 0 0 4224 0 8 6 0 0 4
287 178
368 178
368 194
433 194
2 0 6 0 0 4096 7 8 0 0 7 2
253 174
226 174
0 2 6 0 0 4224 7 0 7 11 0 3
226 111
226 292
345 292
3 0 9 0 0 4096 2 8 0 0 10 2
253 182
201 182
3 0 9 0 0 4096 2 7 0 0 10 2
345 300
201 300
3 1 9 0 0 8320 2 9 5 0 0 3
344 123
201 123
201 344
2 1 6 0 0 0 7 9 4 0 0 3
344 115
226 115
226 83
1 5 9 0 0 4224 8 7 6 0 0 3
379 296
457 296
457 236
1 1 9 0 0 4224 0 9 6 0 0 3
378 119
457 119
457 173
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
196938 1079360 100 100 0 0
0 0 0 0
1 66 162 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 2 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
