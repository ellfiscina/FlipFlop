CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
177209362 0
0
6 Title:
5 Name:
0
0
0
26
13 Logic Switch~
5 224 526 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-5 -17 9 -9
3 V12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3820 0 0
2
41827.9 0
0
13 Logic Switch~
5 223 441 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7678 0 0
2
41827.9 0
0
13 Logic Switch~
5 368 527 0 1 11
0 12
0
0 0 21360 90
2 0V
14 0 28 8
3 V10
10 -10 31 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
961 0 0
2
41827.9 0
0
13 Logic Switch~
5 267 526 0 1 11
0 17
0
0 0 21360 90
2 0V
11 0 25 8
2 V9
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3178 0 0
2
41827.9 0
0
13 Logic Switch~
5 369 435 0 1 11
0 13
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V8
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3409 0 0
2
41827.9 0
0
13 Logic Switch~
5 268 438 0 1 11
0 18
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V7
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3951 0 0
2
41827.9 0
0
13 Logic Switch~
5 317 314 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8885 0 0
2
41827.9 0
0
13 Logic Switch~
5 317 114 0 1 11
0 20
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3780 0 0
2
41827.9 0
0
13 Logic Switch~
5 441 316 0 1 11
0 22
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9265 0 0
2
41827.9 0
0
13 Logic Switch~
5 452 108 0 1 11
0 23
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9442 0 0
2
41827.8 0
0
10 2-In NAND~
219 738 257 0 3 22
0 3 4 2
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
9424 0 0
2
41827.9 0
0
10 2-In NAND~
219 735 163 0 3 22
0 5 2 3
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
9968 0 0
2
41827.9 0
0
10 2-In NAND~
219 635 266 0 3 22
0 6 25 4
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
9281 0 0
2
41827.9 0
0
10 2-In NAND~
219 633 154 0 3 22
0 24 6 5
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
8464 0 0
2
41827.9 0
0
14 Logic Display~
6 478 484 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7168 0 0
2
41827.9 0
0
14 Logic Display~
6 445 449 0 1 2
12 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3171 0 0
2
41827.9 0
0
5 4027~
219 369 507 0 7 32
0 13 10 11 9 12 7 8
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U5B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 2 5 0
1 U
4139 0 0
2
41827.9 0
0
5 4027~
219 268 507 0 7 32
0 18 16 14 15 17 9 10
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U5A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 5 0
1 U
6435 0 0
2
41827.9 0
0
7 Pulser~
4 120 489 0 10 12
0 28 29 14 11 0 0 5 5 3
8
0
0 0 4656 0
0
2 V6
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
5283 0 0
2
41827.9 0
0
7 Pulser~
4 136 205 0 10 12
0 30 31 21 6 0 0 5 5 3
8
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
6874 0 0
2
41827.9 0
0
5 4023~
219 373 275 0 4 22
0 3 21 19 26
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U3A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 1 3 0
1 U
5305 0 0
2
41827.8 0
0
5 4023~
219 373 145 0 4 22
0 20 21 2 27
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U2C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 3 2 0
1 U
34 0 0
2
41827.8 0
0
5 4023~
219 520 275 0 4 22
0 24 26 22 25
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 2 2 0
1 U
969 0 0
2
41827.8 0
0
5 4023~
219 509 145 0 4 22
0 23 27 25 24
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 1 2 0
1 U
8402 0 0
2
41827.8 0
0
14 Logic Display~
6 841 216 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Qn
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3751 0 0
2
41827.8 4
0
14 Logic Display~
6 841 119 0 1 2
12 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 Q
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4292 0 0
2
41827.8 5
0
38
3 0 2 0 0 0 0 11 0 0 37 2
765 257
765 257
3 0 3 0 0 0 0 12 0 0 38 2
762 163
762 163
3 0 4 0 0 0 0 13 0 0 33 2
662 266
662 266
3 0 5 0 0 0 0 14 0 0 34 2
660 154
660 154
0 1 6 0 0 4112 0 0 13 6 0 3
598 205
598 257
611 257
4 2 6 0 0 4224 0 20 14 0 0 4
166 205
598 205
598 163
609 163
6 1 7 0 0 4224 0 17 15 0 0 5
399 489
455 489
455 510
478 510
478 502
7 1 8 0 0 4224 0 17 16 0 0 3
393 471
445 471
445 467
6 4 9 0 0 4224 0 18 17 0 0 2
298 489
345 489
7 2 10 0 0 4224 0 18 17 0 0 2
292 471
345 471
4 3 11 0 0 12416 0 19 17 0 0 6
150 489
189 489
189 554
331 554
331 480
345 480
1 5 12 0 0 4224 0 3 17 0 0 2
369 514
369 513
1 1 13 0 0 4224 0 5 17 0 0 2
369 447
369 450
3 3 14 0 0 4224 0 18 19 0 0 2
244 480
144 480
1 4 15 0 0 8320 0 1 18 0 0 4
236 526
240 526
240 489
244 489
1 2 16 0 0 8320 0 2 18 0 0 4
235 441
240 441
240 471
244 471
1 5 17 0 0 0 0 4 18 0 0 2
268 513
268 513
1 1 18 0 0 0 0 6 18 0 0 2
268 450
268 450
1 3 19 0 0 8320 0 7 21 0 0 4
329 314
339 314
339 284
349 284
1 1 20 0 0 8320 0 8 22 0 0 4
329 114
340 114
340 136
349 136
0 2 21 0 0 8320 0 0 22 22 0 3
248 196
248 145
349 145
3 2 21 0 0 0 0 20 21 0 0 4
160 196
248 196
248 275
349 275
1 3 22 0 0 8320 0 9 23 0 0 4
453 316
464 316
464 284
496 284
1 1 23 0 0 4224 0 10 24 0 0 3
464 108
464 136
485 136
0 1 3 0 0 4224 0 0 21 35 0 4
699 191
326 191
326 266
349 266
0 3 2 0 0 4224 0 0 22 36 0 4
686 224
338 224
338 154
349 154
1 0 24 0 0 8320 0 23 0 0 32 5
496 266
476 266
476 167
574 167
574 145
3 0 25 0 0 12416 0 24 0 0 31 5
485 154
464 154
464 245
574 245
574 275
4 2 26 0 0 4224 0 21 23 0 0 2
400 275
496 275
4 2 27 0 0 4224 0 22 24 0 0 2
400 145
485 145
4 2 25 0 0 0 0 23 13 0 0 2
547 275
611 275
4 1 24 0 0 0 0 24 14 0 0 2
536 145
609 145
0 2 4 0 0 4224 0 0 11 0 0 2
659 266
714 266
0 1 5 0 0 4224 0 0 12 0 0 2
656 154
711 154
1 0 3 0 0 0 0 11 0 0 38 5
714 248
699 248
699 191
794 191
794 163
0 2 2 0 0 0 0 0 12 37 0 5
794 257
794 224
686 224
686 172
711 172
0 1 2 0 0 0 0 0 25 0 0 3
762 257
841 257
841 234
0 1 3 0 0 0 0 0 26 0 0 3
758 163
841 163
841 137
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
